library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity lpf is
begin
    port(
        clk : in std_logic;
        )
end entity;
