type coeff_array is array (0 to 62) of integer;
constant filter_coeff : coeff_array := (
    27,
    20,
    4,
    -19,
    -42,
    -53,
    -41,
    0,
    62,
    118,
    136,
    88,
    -27,
    -174,
    -286,
    -292,
    -150,
    118,
    417,
    608,
    558,
    211,
    -364,
    -967,
    -1313,
    -1127,
    -256,
    1255,
    3143,
    4988,
    6332,
    6823,
    6332,
    4988,
    3143,
    1255,
    -256,
    -1127,
    -1313,
    -967,
    -364,
    211,
    558,
    608,
    417,
    118,
    -150,
    -292,
    -286,
    -174,
    -27,
    88,
    136,
    118,
    62,
    0,
    -41,
    -53,
    -42,
    -19,
    4,
    20,
    27);
